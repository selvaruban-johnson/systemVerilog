module test_reg ();
reg [1:0]a;
reg b[1:0];
reg [1:0]c[2:0];
reg [1:0]d[2:0][3:0];
reg [3:0][1:0]e[2:0];
reg [1:0][2:0]f[3:0][4:0];
endmodule