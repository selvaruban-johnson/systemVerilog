class packet;
rand bit [2:0]a,b;
bit [2:0]s;
bit c;
endclass