class packet;
 
 rand bit we;
 rand bit [7:0] data_in;
 rand bit [2:0] address;
 bit [7:0] data_out;

endclass
