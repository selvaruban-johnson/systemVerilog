class packet;
rand bit [7:0]a,b;
bit [15:0]pro;
endclass 