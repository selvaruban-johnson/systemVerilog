class classtest ;
	int i=43;
	task disp();
		$display("i=%d",i);
	endtask
endclass
		