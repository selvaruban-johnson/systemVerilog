module test_short();
shortint k;
initial
begin
	k = 300*300;
	$display ("k = %d",k);
end
endmodule
