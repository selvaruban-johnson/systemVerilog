//interface 
interface intf();
bit [3:0]a,b,sum;
bit [2:0]s;
bit co;
endinterface 