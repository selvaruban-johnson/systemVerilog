module square_of_3bit (input [2:0]a,output logic [5:0]square);
assign square = a*a;
endmodule 