interface intf ();
bit [7:0]a,b;
bit [15:0]pro;
endinterface 