/*3. Define a class with variable a with size of 3. Randomize class 8 times such that each time a
holds a different value.*/

class class_d10_3;

randc reg [5:0] a;


endclass
