/*1. Define a class with variable a and b and generate random value 5 times and print them.
Overwrite the value of a to 55 after randomization.*/


class class_d10;

int a,b;
task disp();
	$display ("a=%d,b=%d",a,b);
endtask
endclass
