/*2. Define a class with variable u, v and w and generate random value of u and v with fix value of
w (=70).*/

class class_d10_2;

int u,v,w=70;
task disp();
	$display("u=%d v=%d w=%d",u,v,w);
endtask
endclass

