module test_design
(input a,b,c,d,e,f,g,
output logic y);
assign  y = a&b&c&d&e&f&g;

endmodule 