//packet
class packet;
parameter n=4;
rand bit [n-1:0]a,b;
rand bit [2:0]s;
bit [n-1:0]sum;
bit co;
endclass 