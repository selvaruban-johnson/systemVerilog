/*6. Define a class with dynamic array a. Randomize class such that each element of dynamic array
a has value greater than 7
*/


class class_dynamic_d10_6 ;

rand	int a[];
endclass 