interface ri_interface(input bit clk,we);
bit [2:0]addr;
bit [15:0]d_in;
bit [15:0]d_out;
endinterface 