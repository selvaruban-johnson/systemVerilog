class env_packet;
rand bit [2:0]addr;
rand bit [15:0]d_in;
bit [15:0]d_out;
endclass 