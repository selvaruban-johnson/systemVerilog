module new_new();
int f[5]='{1,2,3,4,5};
int d[]='{10,2,30,40,50};
int a[*]='{1:11,2:22,3:33,4:44,5:55};
int q[$]='{1,3,5,7,9};
initial begin
$display("sum=%d",f.sum);
$display("sum%d",d.sum);
$display("sum=%d",a.sum);
$display("sum=%d",q.sum);
$display("product=%d",f.product);
$display("product=%d",d.product);
$display("product%d",a.product);
$display("product%d",q.product);
$display("and=%d",f.and);
$display("and=%d",d.and);
$display("and=%d",a.and);
$display("and=%d",q.and);
$display("or=%d",f.or);
$display("or=%d",d.or);
$display("or=%d",a.or);
$display("or=%d",q.or);
$display("xor=%d",f.xor);
$display("xor=%d",d.xor);
$display("xor=%d",a.xor);
$display("xor=%d",q.xor);
f.sort();
$display("sort=%p",f);
d.sort();
$display("sort=%p",d);
//$display("%d",a.sort);
q.sort();
$display("sort=%p",q);
f.rsort();
$display("rsort=%p",f);
d.rsort();
$display("rsort=%p",d);
//$display("%d",a.rsort);
q.rsort();
$display("rsort=%p",q);
f.reverse();
$display("reverse=%p",f);
d.reverse();
$display("reverse=%p",d);
//$display("%d",a.reverse);
q.reverse();
$display("reverse=%p",q);
f.shuffle();
$display("shuffle=%p",f);
d.shuffle();
$display("shuffle=%p",d);
//$display("%d",a.shuffle);
q.shuffle();
$display("shuffle=%p",q);
$display("unique=%p",f.unique);
$display("unique=%p",d.unique);
$display("unique=%p",a.unique);
$display("unique=%p",q.unique);
$display("max=%p",f.max);
$display("max=%p",d.max);
$display("max=%p",a.max);
$display("max=%p",q.max);
$display("min=%p",f.min);
$display("min=%p",d.min);
$display("min=%p",a.min);
$display("min=%p",q.min);
end
endmodule
